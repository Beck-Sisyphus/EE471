// EE 471 Lab 1,  Beck Pang, Spring 2015
// Main function for calling different counter onto the board
// @require: only call one counter a time
module DE1_SoC_SRAM_test (CLOCK_50, LEDR, SW, KEY);
	input CLOCK_50;  // connect to system 50 MHz clock
	output reg [9:0] LEDR;
	input [9:0] SW;
	input [3:0] KEY;
	
	wire clk;
	wire [15:0] data;
	reg [6:0] hold;
	reg WrEn;
	reg [10:0] adx;
	reg [15:0] store;
	wire clkControl, autoEnter, rst, slowClk;
	//reg [15:0] data;
	//assign data[6:0] = SW[6:0]
	assign clkControl = SW[7];
	assign autoEnter = SW[8];
	assign rst = SW[9];
	assign data = WrEn ? 16'bZ : store;
	
	SRAM2Kby16 memory(clk, adx,  WrEn, data);
	clkSlower counter(slowClk, CLOCK_50, rst);
	
	always @(posedge clk) begin
		if(rst) begin
			hold = 0;
			adx = 0;
			WrEn = 1;
			LEDR = 0;
		end else if(autoEnter) begin
			WrEn = 0;
			adx = hold;
			store = 7'b1111111 - hold;
			LEDR[6:0] = hold;
			hold = hold + 1'b1;	
		end else begin
			WrEn = 1;
			adx = SW[6:0];
			LEDR[6:0] = data[6:0];
		end
	end
	

	assign clk = clkControl ? slowClk : CLOCK_50;
	
endmodule 

module SendP2SBufferTestbench();
	reg CLOCK_50;  // connect to system 50 MHz clock
	wire [9:0] LEDR;
	reg [9:0] SW;
	reg [3:0] KEY;
	DE1_SoC dut (CLOCK_50, LEDR, SW, KEY);
	// Set up the clocking
	
	parameter d = 20;
	initial begin
		CLOCK_50 = 1;
		SW = 12;
		KEY = 0;
	end
	
	always #(d/2) CLOCK_50 = ~CLOCK_50;
	

	// Set up the inputs to the design
	initial begin
		#(d*10); SW[9] = 1;
		#d; SW[9] = 0; SW[8] = 1;
		#(d*500); SW[8] = 0;
		#d SW[5:0] = 64;
		#d SW[5:0] = 32;
		#d SW[5:0] = 16;
		#d SW[5:0] = 8;
		#d SW[5:0] = 120;
		$stop;
	end
endmodule 