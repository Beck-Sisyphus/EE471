module orGate (busOR,  busA, busB);
	output [31:0] busOR;
	input  [31:0] busA, busB;

endmodule