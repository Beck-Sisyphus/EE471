module subtract (busSUB, busA, busB, zSUB, oSUB, cSUB, nSUB);
	output [31:0] busSUB;
	input  [31:0] busA, busB;
	output zSUB, oSUB, cSUB, nSUB;

endmodule