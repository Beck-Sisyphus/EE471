module loader(clk, rst, loadEnable, IMR, instr2load, loadAdx)
	input clk, rst, loadEnable;
	output IMR;
	output [31:0] instr2load;
	output [6:0] loadAdx;
	
	
endmodule
	