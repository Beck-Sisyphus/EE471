// andorTop0.v
`include "andOr0.v"

module testBench ();

	// connext the two modules
	wire [1:0] X, Y;
	wire [1:0] XandY, XorY;

	// declare an instance of the AND module
	AndOr myAndOr (XandY[1:0], XorY[1:0], X[1:0], Y[1:0]);

	Tester aTester (X[1:0], Y[1:0], XandY[1:0], XorY[1:0]);

	// file for gtkwave

	initial
	begin
		$dumpfile("andOr0.vcd");
		$dumpvars(1, myAndOr);
	end

endmodule

module Tester (
	output reg [1:0] xOut, yOut,   
	input [1:0] XandYin, XorYin // Clock Enable
);
//	reg [1:0] xOut, yOut;

	parameter stimDelay = 20;

	initial // Response
	begin
		$display("\t\t xOut yOut \t XandYin XorYin \t   Time ");
		$monitor("\t\t %b\t %b \t %b \t %b", xOut, yOut, XandYin, XorYin, $time);
	end

	initial // Stimulus
	begin
					xOut = 'b00; yOut = 'b10;
		#stimDelay	xOut = 'b10;
		#stimDelay  yOut = 'b01;
		#stimDelay  xOut = 'b11;

		#(2*stimDelay);
		$finish;
	end

endmodule