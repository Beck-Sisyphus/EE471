module setLT (busSLT, busA, busB);
	output [31:0] busSLT;
	input  [31:0] busA, busB;
	
endmodule