module andGate (busAND, busA, busB);
	output [31:0] busAND;
	input  [31:0] busA, busB;

endmodule