module shiftll (busSLL, busA, busB);
	output [31:0] busSLL;
	input  [31:0] busA, busB;
endmodule