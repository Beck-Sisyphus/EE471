module 2Kx16_SRAM(adx,chpSel,OutEn,WrEn,DataIn,DataOut);
input [11:0] adx;
input chpSel;
input OutEn;
input WrEn;
input [15:0] DataIn;
output [15:0] DataOut;









endmodule
